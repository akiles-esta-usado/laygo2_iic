magic
tech sky130A
timestamp 1658356910
<< checkpaint >>
rect -650 -660 938 1668
<< metal1 >>
rect 57 844 87 1028
rect 201 844 231 1028
rect 57 -20 87 164
rect 201 -20 231 164
<< metal2 >>
rect -20 978 308 1038
rect 54 777 234 807
rect 54 633 234 663
rect 54 345 234 375
rect 54 201 234 231
rect -20 -30 308 30
<< metal3 >>
rect 57 345 87 663
rect 129 201 159 807
use nmos13_fast_boundary  MN0_IBNDL0 skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN0_IBNDR0
timestamp 1655824928
transform 1 0 216 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN0_IM0 skywater130_microtemplates_dense
timestamp 1654175211
transform 1 0 72 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN0_IVD0 skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 144 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN0_IVG0
timestamp 1647525606
transform 1 0 144 0 1 360
box -16 -16 16 16
use via_M1_M2_1  MN0_IVTIED0 skywater130_microtemplates_dense
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 72 0 1 0
box -16 -16 16 16
use pmos13_fast_boundary  MP0_IBNDL0 skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 0 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP0_IBNDR0
timestamp 1655825313
transform 1 0 216 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP0_IM0 skywater130_microtemplates_dense
timestamp 1654091791
transform 1 0 72 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP0_IVD0
timestamp 1647525606
transform 1 0 144 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP0_IVG0
timestamp 1647525606
transform 1 0 144 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP0_IVTIED0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 72 0 -1 1008
box -16 -16 16 16
use via_M2_M3_0  NoName_1 skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 72 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 72 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 144 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_7
timestamp 1647525786
transform 1 0 144 0 1 792
box -19 -19 19 19
<< labels >>
flabel metal3 144 504 144 504 0 FreeSans 240 90 0 0 O:
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 I
flabel metal2 144 0 144 0 0 FreeSans 480 0 0 0 VSS
flabel metal2 144 1008 144 1008 0 FreeSans 480 0 0 0 VDD
<< end >>
